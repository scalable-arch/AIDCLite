`define AIDC_LITE_VERSION_MAJOR 8'h01
`define AIDC_LITE_VERSION_MINOR 8'h01
`define AIDC_LITE_VERSION_MICRO 16'h01
`define AIDC_LITE_GIT_HASH      32'h00000000
