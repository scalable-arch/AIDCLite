class transaction;
    bit [63:0] data [16];
    bit [31:0] addr;
endclass
